`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:59:25 09/28/2016 
// Design Name: 
// Module Name:    Behavioral_S4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Behavioral_S4(
    input [63:0] A,
    input [63:0] B,
    output [63:0] SUM
    );
assign SUM= A+B;

endmodule
