`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:32:04 09/25/2016 
// Design Name: 
// Module Name:    SIXTY_4_CLA 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SIXTY_4_CLA(
	 input [63:0] A,
    input [63:0] B,
    output [64:0] SUM,
	 output CARRY,
	 wire CIN
    );
	
	//CLA_2B s1 ( .A (A[0]), .B 

endmodule
